/* verilator lint_off UNUSEDSIGNAL */

module toplevel (
input               clk     , // Top level system clock input.
input               sw_0    , // Button - for reset
input   wire        uart_rxd, // UART Recieve pin.
output  wire        uart_txd  // UART transmit pin.
);


// Clock frequency in hertz.
parameter CLK_HZ = 2000000;
parameter BIT_RATE =   9600;
parameter PAYLOAD_BITS = 8;

wire [PAYLOAD_BITS-1:0]  uart_rx_data;
wire        uart_rx_valid;
wire        uart_rx_break;

wire        uart_tx_busy;
wire [PAYLOAD_BITS-1:0]  uart_tx_data;
wire        uart_tx_en;

wire rst;

reg [31:0] counter;

reg [7:0] data;

assign rst = !sw_0;

always @(posedge clk) begin
  if(counter == CLK_HZ)
    counter <= 0;
  else
    counter <= counter + 1;
  
  if(uart_rx_valid)
    data <= uart_rx_data;
end

// Loopback
assign uart_tx_en = counter == 0;
assign uart_tx_data = data;

/*
puzzle puzzle_ (
  .rst (rst),
  .clk (clk),
  .output_data (uart_tx_data),
  .output_en (uart_tx_en),
  .output_busy (uart_tx_busy),
  .input_data (uart_rx_data),
  .input_valid (uart_rx_valid)
);
*/

// ------------------------------------------------------------------------- 

//
// UART R:X
uart_rx #(
.BIT_RATE(BIT_RATE),
.PAYLOAD_BITS(PAYLOAD_BITS),
.CLK_HZ  (CLK_HZ  )
) i_uart_rx(
.clk          (clk          ), // Top level system clock input.
.resetn       (!rst         ), // Asynchronous active low reset.
.uart_rxd     (uart_rxd     ), // UART Recieve pin.
.uart_rx_en   (1'b1         ), // Recieve enable
.uart_rx_break(uart_rx_break), // Did we get a BREAK message?
.uart_rx_valid(uart_rx_valid), // Valid data recieved and available.
.uart_rx_data (uart_rx_data )  // The recieved data.
);

//
// UART Transmitter module.
//
uart_tx #(
.BIT_RATE(BIT_RATE),
.PAYLOAD_BITS(PAYLOAD_BITS),
.CLK_HZ  (CLK_HZ  )
) i_uart_tx(
.clk          (clk          ),
.resetn       (sw_0         ),
.uart_txd     (uart_txd     ),
.uart_tx_en   (uart_tx_en   ),
.uart_tx_busy (uart_tx_busy ),
.uart_tx_data (uart_tx_data ) 
);


endmodule
